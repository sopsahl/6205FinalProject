`timescale 1ns / 1ps
`default_nettype none



`default_nettype wire