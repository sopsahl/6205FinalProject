package alu_constants;

  parameter logic [3:0] ALU_ADD  = 4'b0000;
  parameter logic [3:0] ALU_SUB  = 4'b0001;
  parameter logic [3:0] ALU_AND  = 4'b0010;
  parameter logic [3:0] ALU_OR   = 4'b0011;
  parameter logic [3:0] ALU_XOR  = 4'b0100;
  parameter logic [3:0] ALU_SLL  = 4'b0101;
  parameter logic [3:0] ALU_SRL  = 4'b0110;
  parameter logic [3:0] ALU_SRA  = 4'b0111;
  parameter logic [3:0] ALU_SLT  = 4'b1000;

endpackage